module led_display(rst, clk, leds, activate);
	input clk, rst;
	input activate;
	
	output [15:0] leds;
	reg [15:0] leds;
	
	integer cnt;

	always @(posedge clk) begin
		if (~rst) begin
			leds = 16'b0;
			cnt = 0;
		end else begin
			if (~activate) leds = 16'b0;
			else begin
				case (cnt)
					0 : leds = 16'b0000000000000001;
					1 : leds = 16'b0000000000000010;
					2 : leds = 16'b0000000000000100;
					3 : leds = 16'b0000000000001000;
					4 : leds = 16'b0000000000010000;
					5 : leds = 16'b0000000000100000;
					6 : leds = 16'b0000000001000000;
					7 : leds = 16'b0000000010000000;
					8 : leds = 16'b1000000000000000;
					9 : leds = 16'b0100000000000000;
					10: leds = 16'b0010000000000000;
					11: leds = 16'b0001000000000000;
					12: leds = 16'b0000100000000000;
					13: leds = 16'b0000010000000000;
					14: leds = 16'b0000001000000000;
					15: leds = 16'b0000000100000000;
					16: leds = 16'b0000000000000001;
					17: leds = 16'b0000000000000010;
					18: leds = 16'b0000000000000100;
					19: leds = 16'b0000000000001000;
					20: leds = 16'b0000000000010000;
					21: leds = 16'b0000000000100000;
					22: leds = 16'b0000000001000000;
					23: leds = 16'b0000000010000000;
					24: leds = 16'b1000000000000000;
					25: leds = 16'b0100000000000000;
					26: leds = 16'b0010000000000000;
					27: leds = 16'b0001000000000000;
					28: leds = 16'b0000100000000000;
					29: leds = 16'b0000010000000000;
					30: leds = 16'b0000001000000000;
					31: leds = 16'b0000000100000000;
					32: leds = 16'b1000000000000001;
					33: leds = 16'b0100000000000010;
					34: leds = 16'b0010000000000100;
					35: leds = 16'b0001000000001000;
					36: leds = 16'b0000100000010000;
					37: leds = 16'b0000010000100000;
					38: leds = 16'b0000001001000000;
					39: leds = 16'b0000000110000000;
					40: leds = 16'b0000000110000000;
					41: leds = 16'b0000001001000000;
					42: leds = 16'b0000010000100000;
					43: leds = 16'b0000100000010000;
					44: leds = 16'b0001000000001000;
					45: leds = 16'b0010000000000100;
					46: leds = 16'b0100000000000010;
					47: leds = 16'b1000000000000001;
				endcase

				if (cnt == 47) cnt = 0;
				else cnt = cnt + 1;
			end
		end
	end
endmodule
